library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.numeric_std.unsigned;
use std.textio.all;

entity div16_8_8 is
	generic(
		A_WIDTH			: POSITIVE := 17;
		B_WIDTH			: POSITIVE := 8;
		RESULT_WIDTH	: POSITIVE := 9
	);
	port (
		clk        : in  STD_LOGIC;
		en         : in  STD_LOGIC;
		rstn       : in  STD_LOGIC;
		a          : in  STD_LOGIC_VECTOR( A_WIDTH-1 downto 0);
		b          : in  STD_LOGIC_VECTOR( B_WIDTH-1 downto 0);
		result     : out STD_LOGIC_VECTOR( RESULT_WIDTH-1 downto 0)		
	);
end entity div16_8_8;

architecture rtl of div16_8_8 is

    type unsigned_8_array  is array(natural range <>) of UNSIGNED( 7 downto 0);
	type unsigned_16_array is array(natural range <>) of UNSIGNED(15 downto 0);

	signal r_remainder 		: unsigned_16_array(1 to 9);
	signal r_shifted_b 		: unsigned_16_array(1 to 9);
	signal r_result    		: unsigned_8_array (1 to 9);
	signal r_result_signed 	: SIGNED(8 downto 0);
	signal r_sign      		: STD_LOGIC_VECTOR(1 to 9);
	signal r_en		     	: STD_LOGIC_VECTOR(1 to 9);
begin

	process(clk, rstn, en)
		variable v_result 	: UNSIGNED( 8 downto 1);
        variable a_signed 	: SIGNED(16 downto 0);
        variable a_unsigned : UNSIGNED(15 downto 0);


	begin
		if rstn = '0' then
	
	        -- STUDENT CODE HERE
			result <= (others => '0');
			r_en <= (others => '0');

			FOR i IN 1 TO 9 LOOP
				r_remainder(i) <= (others => '0');
				r_shifted_b(i) <= (others => '0');
				r_result(i) <= (others => '0');


			END LOOP;

            -- STUDENT CODE until HERE
		elsif rising_edge(clk) and en = '1' then
		
    		-- STUDENT CODE HERE
			-- Initialisieren
				r_remainder(1) 	<= (others => '0');
				r_shifted_b(1) 	<= (others => '0');
				r_result(1) 	<= (others => '0');

			-- Reinschaufeln
				r_remainder(1) <= unsigned(a(15 downto 0));
				r_shifted_b(1)(15 downto 8) <= unsigned(b);
				r_en(1) <= '1';

			-- Berechnen
				-- Vergleicher

				FOR i IN 1 TO 8 LOOP
					IF r_en(i) = '1' THEN
						IF r_remainder(i) <  r_shifted_b(i) THEN
							r_result(i)(8 - i) <= '0';
							r_remainder(i + 1) <= r_remainder(i);
						ELSE
							r_result(i)(8 - i) <= '1';
							r_remainder(i + 1) <= r_remainder(i) - r_shifted_b(i);

						END IF;
					END IF;
				END LOOP;

				r_en(2 to 9) <= r_en(1 to 8);

				-- Shift Divisor
				FOR i IN 1 to 8 LOOP
					r_shifted_b(i + 1) <= (others => '0');
					r_shifted_b(i + 1)((15 - i) downto (8 - i)) <= r_shifted_b(i)((16 - i) downto (9 - i));
				END LOOP;

			
			-- Weitergeben
			--r_remainder(2 to 9) <= r_remainder(1 to 8);
			r_result(2 to 9) <= r_result(1 to 8);
	
			-- Rausschaufeln
			--r_result_signed <= '0' & unsigned(r_result(9));
			-- STUDENT CODE until HERE
		end if;
	end process;
	
	result <= STD_LOGIC_VECTOR(r_result_signed);

end architecture rtl;
